module controlador_over_the_rainbow 
( output Clk_out,
  output reg Disparo,
  output reg [27:0] Temp_out,
  output reg [27:0] Freq_out,	
  input	Clk_in, Duracao, Stop_in, Play_in
);

	///clock da placa
	`define clk_FPGA 50000000 //50MHz
	//overflow para frequencias (50MHz)
	`define Re3 27244 //583Hz (Ré3)
	`define Mi3 24279 //659Hz (Mi3)
	`define Fa3 22922 //698Hz (Fá3)
	`define Sol3 20408 //784Hz (Sol3)
	`define La3 18181 //880Hz (Lá3)
	`define Sib3 17167 //932Hz (Sib3)
	`define Do4 15296 //1046Hz (Dó4)
	`define Re4 13617 //1175Hz (Ré4)
	`define Mi4 12139 //1318Hz (Mi4)
	`define Fa4 11453 //1397Hz (Fá4)
	
	// overflow para tempos (50MHz)
	// BPM igual a 60 implica que t1, 1 batida, representa 1 seg
	//`define BPM 100 //batidas por minuto
	//`define BPS <= BPM / 60 //batidas por segundo
	`define ov_t4 (4 * 16000000) / (100/60) //overflow 4 batidas
	`define ov_t2  (2 * 16000000) / (100/60) //overflow 2 batidas
	`define ov_t1 (16000000) / (100/60) //overflow 1 batida
	`define ov_t1_2 (16000000/2) / (100/60) //overflow 1/2 batidas
	
	//FSM Declaração de estados 
	reg [4:0] estado, prox_estado;
	localparam s0 = 5'b00000;   //define estado 0
	localparam s1 = 5'b00001;   //define estado 1
	localparam s2 = 5'b00010;   //define estado 2
	localparam s3 = 5'b00011;   //define estado 3
	localparam s4 = 5'b00100;   //define estado 4
	localparam s5 = 5'b00101;   //define estado 5
	localparam s6 = 5'b00110;   //define estado 6
	localparam s7 = 5'b00111;   //define estado 7
	localparam s8 = 5'b01000;   //define estado 8
	localparam s9 = 5'b01001;   //define estado 9
	localparam s10 = 5'b01010;   //define estado 10
	localparam s11 = 5'b01011;   //define estado 11
	localparam s12 = 5'b01100;   //define estado 12
	localparam s13 = 5'b01101;   //define estado 13
	localparam s14 = 5'b01110;   //define estado 14
	localparam s15 = 5'b01111;   //define estado 15
	localparam s16 = 5'b10000;   //define estado 16
	localparam s17 = 5'b10001;   //define estado 17
	localparam s18 = 5'b10010;   //define estado 18
	localparam s19 = 5'b10011;   //define estado 19
	localparam s20 = 5'b10100;   //define estado 20
	localparam s21 = 5'b10101;   //define estado 21
	localparam s22 = 5'b10110;   //define estado 22
	localparam s23 = 5'b10111;   //define estado 23
	localparam s24 = 5'b11000;   //define estado 24
	
	always @ (posedge Clk_in)
	begin : L1
		estado <= prox_estado;
	end
	
	always @ (*)//Combinacional 
	begin : L2
		case (estado)
			s0: if (Stop_in == 1'b1)
				 begin
					prox_estado <= s0;
				 end
				 else
				 begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s1;
					else prox_estado <= s0;
				end
			s1: if (Stop_in == 1'b1)
				 begin
					prox_estado <= s0;
				 end
				 else
				 begin 
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s2;
					else prox_estado <= s1;
				 end
			s2: if (Stop_in == 1'b1)
				 begin
					prox_estado <= s0;
				 end
				 else
				 begin
					if (Duracao == 1'b0 && Play_in == 1'b1) 
						prox_estado <= s3;
					else prox_estado <= s2;
				 end
			s3:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1) 
						prox_estado <= s4;
					else prox_estado <= s3;
				end
			s4:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s5;
					else prox_estado <= s4;
				end
			s5:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1) 
						prox_estado <= s6;
					else prox_estado <= s5;
				end
			s6:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1) 
						prox_estado <= s7;
					else prox_estado <= s6;
				end
			s7:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1) 
						prox_estado <= s8;
					else prox_estado <= s7;
				end
			s8:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end 
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s9;
					else prox_estado <= s8;
				end
			s9:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s10;
					else prox_estado <= s9;
				end
			s10:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s11;
					else prox_estado <= s10;
				end
			s11:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s12;
					else prox_estado <= s11;
				end
			s12:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s13;
					else prox_estado <= s12;
				end
			s13:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s14;
					else prox_estado <= s13;
				end
			s14:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s15;
					else prox_estado <= s14;
				end
			s15:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end 
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s16;
					else prox_estado <= s15;
				end
			s16:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s17;
					else prox_estado <= s16;
				end
			s17:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s18;
					else prox_estado <= s17;
				end
			s18:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end 
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s19;
					else prox_estado <= s18;
				end
			s19:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s20;
					else prox_estado <= s19;
				end
			s20:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end 
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s21;
					else prox_estado <= s20;
				end
			s21:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end 
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s22;
					else prox_estado <= s21;
				end
			s22:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s23;
					else prox_estado <= s22;
				end
			s23:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s24;
					else prox_estado <= s23;
				end
			s24:if (Stop_in == 1'b1)
				begin
					prox_estado <= s0;
				end
				else
				begin
					if (Duracao == 1'b0 && Play_in == 1'b1)
						prox_estado <= s1;
					else prox_estado <= s24;
				end
			default: prox_estado <= s0; //recupera de estado inválido
		endcase
	end	
	
	//FSM Lógica para controle das saídas
	always @ (estado)//Combinacional 
	begin : L3
		case (estado) //s0 apenas inicia a prox nota
			s0: nota(0,`ov_t1);  //freq atual, dur prox		
			s1: nota(`Fa3,`ov_t2);//freq atual, dur prox
			s2: nota(`Fa4,`ov_t2);//freq atual, dur prox
			s3: nota(`Mi4,`ov_t1);//freq atual, dur prox
			s4: nota(`Do4,`ov_t1_2);//freq atual, dur prox
			s5: nota(`Re4,`ov_t1_2);//freq atual, dur prox
			s6: nota(`Mi4,`ov_t1);//freq atual, dur prox
			s7: nota(`Fa4,`ov_t1);//freq atual, dur prox
			s8: nota(`Fa3,`ov_t2);//freq atual, dur prox
			s9: nota(`Re4,`ov_t2);//freq atual, dur prox
			s10: nota(`Do4,`ov_t4);//freq atual, dur prox
			s11: nota(`Re3,`ov_t2);//freq atual, dur prox
			s12: nota(`Sib3,`ov_t2);//freq atual, dur prox
			s13: nota(`La3,`ov_t1);//freq atual, dur prox
			s14: nota(`Fa3,`ov_t1_2);//freq atual, dur prox
			s15: nota(`Sol3,`ov_t1_2);//freq atual, dur prox
			s16: nota(`La3,`ov_t1);//freq atual, dur prox
			s17: nota(`Sib3,`ov_t1);//freq atual, dur prox
			s18: nota(`Sol3,`ov_t1);//freq atual, dur prox
			s19: nota(`Mi3,`ov_t1_2);//freq atual, dur prox
			s20: nota(`Fa3,`ov_t1_2);//freq atual, dur prox
			s21: nota(`Sol3,`ov_t1);//freq atual, dur prox
			s22: nota(`La3,`ov_t1);//freq atual, dur prox
			s23: nota(`Fa3,`ov_t4);//freq atual, dur prox
			s24: nota(0,`ov_t4);//freq atual, dur prox
		endcase
	end
	
	
	//Atribuição contínua
	assign Clk_out = Duracao & Clk_in;	
	
	//Tarefa para atribuição de saídas nos estados
	task nota( input [27:0] ov_f, ov_t);
	begin
		Temp_out = ov_t; //define a duração	proxima nota			
		Freq_out = ov_f; //define a frequência nota atual
		Disparo = 1'b1;  //dispara o temp a próxima nota		
	end
	endtask
	
endmodule		